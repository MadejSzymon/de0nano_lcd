// megafunction wizard: %LPM_MUX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: LPM_MUX 

// ============================================================
// File Name: data_mux.v
// Megafunction Name(s):
// 			LPM_MUX
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 18.1.0 Build 625 09/12/2018 SJ Lite Edition
// ************************************************************


//Copyright (C) 2018  Intel Corporation. All rights reserved.
//Your use of Intel Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Intel Program License 
//Subscription Agreement, the Intel Quartus Prime License Agreement,
//the Intel FPGA IP License Agreement, or other applicable license
//agreement, including, without limitation, that your use is for
//the sole purpose of programming logic devices manufactured by
//Intel and sold by Intel or its authorized distributors.  Please
//refer to the applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module data_mux (
	clock,
	data0x,
	data10x,
	data11x,
	data12x,
	data13x,
	data14x,
	data15x,
	data16x,
	data17x,
	data18x,
	data19x,
	data1x,
	data20x,
	data21x,
	data22x,
	data23x,
	data24x,
	data25x,
	data26x,
	data27x,
	data28x,
	data29x,
	data2x,
	data30x,
	data31x,
	data32x,
	data33x,
	data34x,
	data35x,
	data36x,
	data37x,
	data38x,
	data39x,
	data3x,
	data4x,
	data5x,
	data6x,
	data7x,
	data8x,
	data9x,
	sel,
	result);

	input	  clock;
	input	[8:0]  data0x;
	input	[8:0]  data10x;
	input	[8:0]  data11x;
	input	[8:0]  data12x;
	input	[8:0]  data13x;
	input	[8:0]  data14x;
	input	[8:0]  data15x;
	input	[8:0]  data16x;
	input	[8:0]  data17x;
	input	[8:0]  data18x;
	input	[8:0]  data19x;
	input	[8:0]  data1x;
	input	[8:0]  data20x;
	input	[8:0]  data21x;
	input	[8:0]  data22x;
	input	[8:0]  data23x;
	input	[8:0]  data24x;
	input	[8:0]  data25x;
	input	[8:0]  data26x;
	input	[8:0]  data27x;
	input	[8:0]  data28x;
	input	[8:0]  data29x;
	input	[8:0]  data2x;
	input	[8:0]  data30x;
	input	[8:0]  data31x;
	input	[8:0]  data32x;
	input	[8:0]  data33x;
	input	[8:0]  data34x;
	input	[8:0]  data35x;
	input	[8:0]  data36x;
	input	[8:0]  data37x;
	input	[8:0]  data38x;
	input	[8:0]  data39x;
	input	[8:0]  data3x;
	input	[8:0]  data4x;
	input	[8:0]  data5x;
	input	[8:0]  data6x;
	input	[8:0]  data7x;
	input	[8:0]  data8x;
	input	[8:0]  data9x;
	input	[5:0]  sel;
	output	[8:0]  result;

	wire [8:0] sub_wire41;
	wire [8:0] sub_wire40 = data39x[8:0];
	wire [8:0] sub_wire39 = data38x[8:0];
	wire [8:0] sub_wire38 = data37x[8:0];
	wire [8:0] sub_wire37 = data36x[8:0];
	wire [8:0] sub_wire36 = data35x[8:0];
	wire [8:0] sub_wire35 = data34x[8:0];
	wire [8:0] sub_wire34 = data33x[8:0];
	wire [8:0] sub_wire33 = data32x[8:0];
	wire [8:0] sub_wire32 = data31x[8:0];
	wire [8:0] sub_wire31 = data30x[8:0];
	wire [8:0] sub_wire30 = data29x[8:0];
	wire [8:0] sub_wire29 = data28x[8:0];
	wire [8:0] sub_wire28 = data27x[8:0];
	wire [8:0] sub_wire27 = data26x[8:0];
	wire [8:0] sub_wire26 = data25x[8:0];
	wire [8:0] sub_wire25 = data24x[8:0];
	wire [8:0] sub_wire24 = data23x[8:0];
	wire [8:0] sub_wire23 = data22x[8:0];
	wire [8:0] sub_wire22 = data21x[8:0];
	wire [8:0] sub_wire21 = data20x[8:0];
	wire [8:0] sub_wire20 = data19x[8:0];
	wire [8:0] sub_wire19 = data18x[8:0];
	wire [8:0] sub_wire18 = data17x[8:0];
	wire [8:0] sub_wire17 = data16x[8:0];
	wire [8:0] sub_wire16 = data15x[8:0];
	wire [8:0] sub_wire15 = data14x[8:0];
	wire [8:0] sub_wire14 = data13x[8:0];
	wire [8:0] sub_wire13 = data12x[8:0];
	wire [8:0] sub_wire12 = data11x[8:0];
	wire [8:0] sub_wire11 = data10x[8:0];
	wire [8:0] sub_wire10 = data9x[8:0];
	wire [8:0] sub_wire9 = data8x[8:0];
	wire [8:0] sub_wire8 = data7x[8:0];
	wire [8:0] sub_wire7 = data6x[8:0];
	wire [8:0] sub_wire6 = data5x[8:0];
	wire [8:0] sub_wire5 = data4x[8:0];
	wire [8:0] sub_wire4 = data3x[8:0];
	wire [8:0] sub_wire3 = data2x[8:0];
	wire [8:0] sub_wire2 = data1x[8:0];
	wire [8:0] sub_wire0 = data0x[8:0];
	wire [359:0] sub_wire1 = {sub_wire40, sub_wire39, sub_wire38, sub_wire37, sub_wire36, sub_wire35, sub_wire34, sub_wire33, sub_wire32, sub_wire31, sub_wire30, sub_wire29, sub_wire28, sub_wire27, sub_wire26, sub_wire25, sub_wire24, sub_wire23, sub_wire22, sub_wire21, sub_wire20, sub_wire19, sub_wire18, sub_wire17, sub_wire16, sub_wire15, sub_wire14, sub_wire13, sub_wire12, sub_wire11, sub_wire10, sub_wire9, sub_wire8, sub_wire7, sub_wire6, sub_wire5, sub_wire4, sub_wire3, sub_wire2, sub_wire0};
	wire [8:0] result = sub_wire41[8:0];

	lpm_mux	LPM_MUX_component (
				.clock (clock),
				.data (sub_wire1),
				.sel (sel),
				.result (sub_wire41)
				// synopsys translate_off
				,
				.aclr (),
				.clken ()
				// synopsys translate_on
				);
	defparam
		LPM_MUX_component.lpm_pipeline = 1,
		LPM_MUX_component.lpm_size = 40,
		LPM_MUX_component.lpm_type = "LPM_MUX",
		LPM_MUX_component.lpm_width = 9,
		LPM_MUX_component.lpm_widths = 6;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: new_diagram STRING "1"
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: CONSTANT: LPM_PIPELINE NUMERIC "1"
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "40"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "9"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "6"
// Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
// Retrieval info: USED_PORT: data0x 0 0 9 0 INPUT NODEFVAL "data0x[8..0]"
// Retrieval info: USED_PORT: data10x 0 0 9 0 INPUT NODEFVAL "data10x[8..0]"
// Retrieval info: USED_PORT: data11x 0 0 9 0 INPUT NODEFVAL "data11x[8..0]"
// Retrieval info: USED_PORT: data12x 0 0 9 0 INPUT NODEFVAL "data12x[8..0]"
// Retrieval info: USED_PORT: data13x 0 0 9 0 INPUT NODEFVAL "data13x[8..0]"
// Retrieval info: USED_PORT: data14x 0 0 9 0 INPUT NODEFVAL "data14x[8..0]"
// Retrieval info: USED_PORT: data15x 0 0 9 0 INPUT NODEFVAL "data15x[8..0]"
// Retrieval info: USED_PORT: data16x 0 0 9 0 INPUT NODEFVAL "data16x[8..0]"
// Retrieval info: USED_PORT: data17x 0 0 9 0 INPUT NODEFVAL "data17x[8..0]"
// Retrieval info: USED_PORT: data18x 0 0 9 0 INPUT NODEFVAL "data18x[8..0]"
// Retrieval info: USED_PORT: data19x 0 0 9 0 INPUT NODEFVAL "data19x[8..0]"
// Retrieval info: USED_PORT: data1x 0 0 9 0 INPUT NODEFVAL "data1x[8..0]"
// Retrieval info: USED_PORT: data20x 0 0 9 0 INPUT NODEFVAL "data20x[8..0]"
// Retrieval info: USED_PORT: data21x 0 0 9 0 INPUT NODEFVAL "data21x[8..0]"
// Retrieval info: USED_PORT: data22x 0 0 9 0 INPUT NODEFVAL "data22x[8..0]"
// Retrieval info: USED_PORT: data23x 0 0 9 0 INPUT NODEFVAL "data23x[8..0]"
// Retrieval info: USED_PORT: data24x 0 0 9 0 INPUT NODEFVAL "data24x[8..0]"
// Retrieval info: USED_PORT: data25x 0 0 9 0 INPUT NODEFVAL "data25x[8..0]"
// Retrieval info: USED_PORT: data26x 0 0 9 0 INPUT NODEFVAL "data26x[8..0]"
// Retrieval info: USED_PORT: data27x 0 0 9 0 INPUT NODEFVAL "data27x[8..0]"
// Retrieval info: USED_PORT: data28x 0 0 9 0 INPUT NODEFVAL "data28x[8..0]"
// Retrieval info: USED_PORT: data29x 0 0 9 0 INPUT NODEFVAL "data29x[8..0]"
// Retrieval info: USED_PORT: data2x 0 0 9 0 INPUT NODEFVAL "data2x[8..0]"
// Retrieval info: USED_PORT: data30x 0 0 9 0 INPUT NODEFVAL "data30x[8..0]"
// Retrieval info: USED_PORT: data31x 0 0 9 0 INPUT NODEFVAL "data31x[8..0]"
// Retrieval info: USED_PORT: data32x 0 0 9 0 INPUT NODEFVAL "data32x[8..0]"
// Retrieval info: USED_PORT: data33x 0 0 9 0 INPUT NODEFVAL "data33x[8..0]"
// Retrieval info: USED_PORT: data34x 0 0 9 0 INPUT NODEFVAL "data34x[8..0]"
// Retrieval info: USED_PORT: data35x 0 0 9 0 INPUT NODEFVAL "data35x[8..0]"
// Retrieval info: USED_PORT: data36x 0 0 9 0 INPUT NODEFVAL "data36x[8..0]"
// Retrieval info: USED_PORT: data37x 0 0 9 0 INPUT NODEFVAL "data37x[8..0]"
// Retrieval info: USED_PORT: data38x 0 0 9 0 INPUT NODEFVAL "data38x[8..0]"
// Retrieval info: USED_PORT: data39x 0 0 9 0 INPUT NODEFVAL "data39x[8..0]"
// Retrieval info: USED_PORT: data3x 0 0 9 0 INPUT NODEFVAL "data3x[8..0]"
// Retrieval info: USED_PORT: data4x 0 0 9 0 INPUT NODEFVAL "data4x[8..0]"
// Retrieval info: USED_PORT: data5x 0 0 9 0 INPUT NODEFVAL "data5x[8..0]"
// Retrieval info: USED_PORT: data6x 0 0 9 0 INPUT NODEFVAL "data6x[8..0]"
// Retrieval info: USED_PORT: data7x 0 0 9 0 INPUT NODEFVAL "data7x[8..0]"
// Retrieval info: USED_PORT: data8x 0 0 9 0 INPUT NODEFVAL "data8x[8..0]"
// Retrieval info: USED_PORT: data9x 0 0 9 0 INPUT NODEFVAL "data9x[8..0]"
// Retrieval info: USED_PORT: result 0 0 9 0 OUTPUT NODEFVAL "result[8..0]"
// Retrieval info: USED_PORT: sel 0 0 6 0 INPUT NODEFVAL "sel[5..0]"
// Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 9 0 data0x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 90 data10x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 99 data11x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 108 data12x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 117 data13x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 126 data14x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 135 data15x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 144 data16x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 153 data17x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 162 data18x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 171 data19x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 9 data1x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 180 data20x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 189 data21x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 198 data22x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 207 data23x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 216 data24x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 225 data25x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 234 data26x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 243 data27x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 252 data28x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 261 data29x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 18 data2x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 270 data30x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 279 data31x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 288 data32x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 297 data33x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 306 data34x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 315 data35x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 324 data36x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 333 data37x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 342 data38x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 351 data39x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 27 data3x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 36 data4x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 45 data5x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 54 data6x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 63 data7x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 72 data8x 0 0 9 0
// Retrieval info: CONNECT: @data 0 0 9 81 data9x 0 0 9 0
// Retrieval info: CONNECT: @sel 0 0 6 0 sel 0 0 6 0
// Retrieval info: CONNECT: result 0 0 9 0 @result 0 0 9 0
// Retrieval info: GEN_FILE: TYPE_NORMAL data_mux.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL data_mux.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL data_mux.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL data_mux.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL data_mux_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL data_mux_bb.v FALSE
// Retrieval info: LIB_FILE: lpm
